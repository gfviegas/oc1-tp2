module main;
  initial
    begin
      $display("Teste");
      $finish;
    end
endmodule
