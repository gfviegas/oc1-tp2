module pc (
  input wire [31:0] naoFacoIdeia,
  output wire [31:0] naoSei
);

endmodule
